module sqs(
    input        b_up,
    input  [2:0] p_state,
    output [2:0] m_state
);
