module op_01(
    input a
        )
