module states()


